library ieee;
use ieee.std_logic_1164.all;

entity demuxOP is 
	port(
		OP: in std_logic_vector (3 downto 0);
		slt_op: out std_logic_vector (2 downto 0);
		rc_ops: out std_logic;
		const_ops: out std_logic;
		sln_ops: out std_logic;
		nand_op: out std_logic;
		lw_op: out std_logic;
		sw_op: out std_logic
	);

end;

architecture arcDemuxOP of demuxOP is
	begin
		process(OP) is
		begin
			case(OP) is
				when "0000" => slt_op <= "000";
									rc_ops <= '1';
									const_ops <= '0';
									sln_ops <= '0';
									nand_op <= '0';
									lw_op <= '0';
									sw_op <= '0';
				when "0001" => slt_op <= "000";
									rc_ops <= '0';
									const_ops <= '1';
									sln_ops <= '0';
									nand_op <= '0';
									lw_op <= '0';
									sw_op <= '0';
				when "0010" => slt_op <= "001";
									rc_ops <= '1';
									const_ops <= '0';
									sln_ops <= '0';
									nand_op <= '0';
									lw_op <= '0';
									sw_op <= '0';
				when "0011" => slt_op <= "001";
									rc_ops <= '0';
									const_ops <= '1';
									sln_ops <= '0';
									nand_op <= '0';
									lw_op <= '0';
									sw_op <= '0';
				when "0100" => slt_op <= "010";
									rc_ops <= '1';
									const_ops <= '0';
									sln_ops <= '0';
									nand_op <= '0';
									lw_op <= '0';
									sw_op <= '0';
				when "0101" => slt_op <= "010";
									rc_ops <= '0';
									const_ops <= '0';
									sln_ops <= '1';
									nand_op <= '0';
									lw_op <= '0';
									sw_op <= '0';
				when "0110" => slt_op <= "011";
									rc_ops <= '1';
									const_ops <= '0';
									sln_ops <= '0';
									nand_op <= '0';
									lw_op <= '0';
									sw_op <= '0';
				when "0111" => slt_op <= "011";
									rc_ops <= '0';
									const_ops <= '0';
									sln_ops <= '1';
									nand_op <= '0';
									lw_op <= '0';
									sw_op <= '0';
				when "1000" => slt_op <= "100";
									rc_ops <= '1';
									const_ops <= '0';
									sln_ops <= '0';
									nand_op <= '0';
									lw_op <= '0';
									sw_op <= '0';
				when "1001" => slt_op <= "100";
									rc_ops <= '1';
									const_ops <= '0';
									sln_ops <= '0';
									nand_op <= '1';
									lw_op <= '0';
									sw_op <= '0';
				when "1010" => slt_op <= "101";
									rc_ops <= '1';
									const_ops <= '0';
									sln_ops <= '0';
									nand_op <= '0';
									lw_op <= '0';
									sw_op <= '0';
				when "1011" => slt_op <= "110";
									rc_ops <= '1';
									const_ops <= '0';
									sln_ops <= '0';
									nand_op <= '0';
									lw_op <= '0';
									sw_op <= '0';
				when "1100" => slt_op <= "111";
									rc_ops <= '0';
									const_ops <= '0';
									sln_ops <= '0';
									nand_op <= '0';
									lw_op <= '1';
									sw_op <= '0';
				when "1110" => slt_op <= "111";
									rc_ops <= '1';
									const_ops <= '0';
									sln_ops <= '0';
									nand_op <= '0';
									lw_op <= '0';
									sw_op <= '1';
				when others => slt_op <= "111";
									rc_ops <= '0';
									const_ops <= '0';
									sln_ops <= '0';
									nand_op <= '0';
									lw_op <= '0';
									sw_op <= '0';
			end case;
		end process;			
end arcDemuxOP;